`timescale 1ns/1ns
module tb_logic2048();
    parameter STEP = 20;
    reg [79:0] initial_board;
    reg [1:0] movDir;
    reg clk, rst;
    wire [31:0] random;
    reg [1:0] restrected;
    reg [2:0] restrect_prob;
    wire stuck;
    wire calc_done;
    wire movable;
    wire [79:0] board_after;
    wire [79:0] filledBoard, storedBoard, mergedBoard;
    wire [2:0] state;
    wire random_clk;
    logic2048 trialUnit(.clk(clk), .rst(rst), .calc_done(calc_done), .random(random[22:0]), .initial_board(initial_board), .restrected(restrected), .restrect_prob(restrect_prob), .stuck(stuck), .filledBoard(filledBoard), .storedBoard(storedBoard), .mergedBoard(mergedBoard), .state(state), .random_clk(random_clk));
    xorshift32 rnd(.clk(random_clk), .rst(rst), .res(random));
    initial begin
        $dumpfile("tb_logic2048.vcd");
        $dumpvars(0, tb_logic2048);
        rst = 0;
        initial_board = {5'd3, 5'd4, 5'd5, 5'd6, 5'd7 ,5'd8, 5'd9, 5'd10, 5'd11 ,5'd12, 5'd13, 5'd14, 5'd15, 5'd16};
        restrected = 0;
        restrect_prob = 7;
#STEP   clk = 0;
#STEP   rst = 1;
        toggleClk;
        toggleClk;
        rst = 0;
        toggleClk;
        toggleClk;
        showState;
        showStored;
        toggleClk;
        toggleClk;
        showState;
        showStored;
        toggleClk;
        toggleClk;
        showState;
        showStored;
        toggleClk;
        toggleClk;
        showState;
        showStored;
        toggleClk;
        toggleClk;
        showState;
        showStored;
        toggleClk;
        toggleClk;
        showState;
        showStored;
        toggleClk;
        toggleClk;
        showState;
        showStored;
        toggleClk;
        toggleClk;
        showState;
        showStored;
        toggleClk;
        toggleClk;
        showState;
        showStored;
        toggleClk;
        toggleClk;
        showState;
        showStored;
        toggleClk;
        toggleClk;
        showState;
        showStored;
        toggleClk;
        toggleClk;
        showState;
        showStored;
        toggleClk;
        toggleClk;
        showState;
        showStored;
        toggleClk;
        toggleClk;
        showState;
        showStored;
        toggleClk;
        toggleClk;
        showState;
        showStored;
        toggleClk;
        toggleClk;
        showState;
        showStored;
        toggleClk;
        toggleClk;
        showState;
        showStored;
        toggleClk;
        toggleClk;
        showState;
        showStored;
        toggleClk;
        toggleClk;
        showState;
        showStored;
        toggleClk;
        toggleClk;
        showState;
        showStored;
        toggleClk;
        toggleClk;
        showState;
        showStored;
        toggleClk;
        toggleClk;
        showState;
        showStored;
        toggleClk;
        toggleClk;
        showState;
        showStored;
        toggleClk;
        toggleClk;
        showState;
        showStored;
        toggleClk;
        toggleClk;
        showState;
        showStored;
        toggleClk;
        toggleClk;
        showState;
        showStored;
        toggleClk;
        toggleClk;
        showState;
        showStored;
        toggleClk;
        toggleClk;
        showState;
        showStored;
        toggleClk;
        toggleClk;
        showState;
        showStored;
        toggleClk;
        toggleClk;
        showState;
        showStored;
        toggleClk;
        toggleClk;
        showState;
        showStored;
        toggleClk;
        toggleClk;
        showState;
        showStored;
        toggleClk;
        toggleClk;
        showState;
        showStored;
        toggleClk;
        toggleClk;
        showState;
        showStored;
        toggleClk;
        toggleClk;
        showState;
        showStored;
        toggleClk;
        toggleClk;
        showState;
        showStored;
        toggleClk;
        toggleClk;
        showState;
        showStored;
        toggleClk;
        toggleClk;
        showState;
        showStored;
        toggleClk;
        toggleClk;
        showState;
        showStored;
        toggleClk;
        toggleClk;
        showState;
        showStored;
        toggleClk;
        toggleClk;
        showState;
        showStored;
        toggleClk;
        toggleClk;
        showState;
        showStored;
        toggleClk;
        toggleClk;
        showState;
        showStored;
        toggleClk;
        toggleClk;
        showState;
        showStored;
        toggleClk;
        toggleClk;
        showState;
        showStored;
        toggleClk;
        toggleClk;
        showState;
        showStored;
        toggleClk;
        toggleClk;
        showState;
        showStored;
        toggleClk;
        toggleClk;
        showState;
        showStored;
        toggleClk;
        toggleClk;
        showState;
        showStored;
        toggleClk;
        toggleClk;
        showState;
        showStored;
        toggleClk;
        toggleClk;
        showState;
        showStored;
        toggleClk;
        toggleClk;
        showState;
        showStored;
        $dumpflush;
        $finish;
    end
    task showStored;
        begin
            $display("storedBoard:");
            $display("%d %d %d %d",storedBoard[19:15], storedBoard[14:10], storedBoard[9:5], storedBoard[4:0]);
            $display("%d %d %d %d",storedBoard[39:35], storedBoard[34:30], storedBoard[29:25], storedBoard[24:20]);
            $display("%d %d %d %d",storedBoard[59:55], storedBoard[54:50], storedBoard[49:45], storedBoard[44:40]);
            $display("%d %d %d %d",storedBoard[79:75], storedBoard[74:70], storedBoard[69:65], storedBoard[64:60]);
            $display("stuck:%d", stuck);
            $display("");
        end
    endtask
    task showMerged;
        begin
            $display("mergedBoard:");
            $display("%d %d %d %d",mergedBoard[19:15], mergedBoard[14:10], mergedBoard[9:5], mergedBoard[4:0]);
            $display("%d %d %d %d",mergedBoard[39:35], mergedBoard[34:30], mergedBoard[29:25], mergedBoard[24:20]);
            $display("%d %d %d %d",mergedBoard[59:55], mergedBoard[54:50], mergedBoard[49:45], mergedBoard[44:40]);
            $display("%d %d %d %d",mergedBoard[79:75], mergedBoard[74:70], mergedBoard[69:65], mergedBoard[64:60]);
            $display("stuck:%d", stuck);
            $display("");
        end
    endtask
    task toggleClk;
        begin
#STEP       clk <= ~clk;
        end
    endtask
    task showState;
        begin
            $display("state:%d",state);
        end
    endtask
    always @(posedge calc_done) begin
        showMerged;
    end
endmodule
